`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 16.04.2021 15:30:14
// Design Name: 
// Module Name: tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb();
parameter Total_MCUs = 8;
reg start;
reg [1:Total_MCUs] rst;
reg [7:0] I[1:Total_MCUs];
reg [7:0]M[0:64*Total_MCUs - 1];  // 2 MCUs
reg [7:0]ctr;
reg [19:0] overall_ctr;
reg clk;
reg [1:Total_MCUs] en;
reg [0:13] dc_in[1:Total_MCUs];
reg [0:10] MCU_ctr; // To keep track of present MCU
reg first_MCU, st;
reg [9:0] present_MCU;
wire [0:22] O[1:Total_MCUs];
wire ready[1:Total_MCUs];
wire done[1:Total_MCUs];
wire [0:13] dc_out[1:Total_MCUs];
wire [1:Total_MCUs]Valid_output;

reg [1:Total_MCUs]start_MCU;
reg change;
//wire [0:10] Total_MCUs;
//assign Total_MCUs = 11'd2;

reg [4:0] on_ctr, off_ctr;

initial begin
clk =0;
ctr=0;
overall_ctr <= 0;

M[0] = 8'd180; M[1] = 8'd183; M[2] = 8'd189; M[3] = 8'd194; M[4] = 8'd198; M[5] = 8'd189; M[6] = 8'd192; M[7] = 8'd201; 
M[64] = 8'd191; M[65] = 8'd187; M[66] = 8'd183; M[67] = 8'd218; M[68] = 8'd237; M[69] = 8'd213; M[70] = 8'd197; M[71] = 8'd200; 
M[128] = 8'd190; M[129] = 8'd187; M[130] = 8'd196; M[131] = 8'd241; M[132] = 8'd16; M[133] = 8'd232; M[134] = 8'd194; M[135] = 8'd201; 
M[192] = 8'd191; M[193] = 8'd186; M[194] = 8'd199; M[195] = 8'd250; M[196] = 8'd26; M[197] = 8'd234; M[198] = 8'd198; M[199] = 8'd197; 
M[256] = 8'd195; M[257] = 8'd189; M[258] = 8'd196; M[259] = 8'd232; M[260] = 8'd254; M[261] = 8'd216; M[262] = 8'd196; M[263] = 8'd198; 
M[320] = 8'd207; M[321] = 8'd193; M[322] = 8'd188; M[323] = 8'd198; M[324] = 8'd205; M[325] = 8'd196; M[326] = 8'd186; M[327] = 8'd203; 
M[384] = 8'd213; M[385] = 8'd199; M[386] = 8'd192; M[387] = 8'd187; M[388] = 8'd183; M[389] = 8'd189; M[390] = 8'd193; M[391] = 8'd211; 
M[448] = 8'd215; M[449] = 8'd207; M[450] = 8'd197; M[451] = 8'd196; M[452] = 8'd193; M[453] = 8'd204; M[454] = 8'd206; M[455] = 8'd222; 

M[8] = 8'd180; M[9] = 8'd183; M[10] = 8'd189; M[11] = 8'd194; M[12] = 8'd198; M[13] = 8'd189; M[14] = 8'd192; M[15] = 8'd201; 
M[72] = 8'd191; M[73] = 8'd187; M[74] = 8'd183; M[75] = 8'd218; M[76] = 8'd237; M[77] = 8'd213; M[78] = 8'd197; M[79] = 8'd200; 
M[136] = 8'd190; M[137] = 8'd187; M[138] = 8'd196; M[139] = 8'd241; M[140] = 8'd16; M[141] = 8'd232; M[142] = 8'd194; M[143] = 8'd201; 
M[200] = 8'd191; M[201] = 8'd186; M[202] = 8'd199; M[203] = 8'd250; M[204] = 8'd26; M[205] = 8'd234; M[206] = 8'd198; M[207] = 8'd197; 
M[264] = 8'd195; M[265] = 8'd189; M[266] = 8'd196; M[267] = 8'd232; M[268] = 8'd254; M[269] = 8'd216; M[270] = 8'd196; M[271] = 8'd198; 
M[328] = 8'd207; M[329] = 8'd193; M[330] = 8'd188; M[331] = 8'd198; M[332] = 8'd205; M[333] = 8'd196; M[334] = 8'd186; M[335] = 8'd203; 
M[392] = 8'd213; M[393] = 8'd199; M[394] = 8'd192; M[395] = 8'd187; M[396] = 8'd183; M[397] = 8'd189; M[398] = 8'd193; M[399] = 8'd211; 
M[456] = 8'd215; M[457] = 8'd207; M[458] = 8'd197; M[459] = 8'd196; M[460] = 8'd193; M[461] = 8'd204; M[462] = 8'd206; M[463] = 8'd222; 

M[16] = 8'd180; M[17] = 8'd183; M[18] = 8'd189; M[19] = 8'd194; M[20] = 8'd198; M[21] = 8'd189; M[22] = 8'd192; M[23] = 8'd201; 
M[80] = 8'd191; M[81] = 8'd187; M[82] = 8'd183; M[83] = 8'd218; M[84] = 8'd237; M[85] = 8'd213; M[86] = 8'd197; M[87] = 8'd200; 
M[144] = 8'd190; M[145] = 8'd187; M[146] = 8'd196; M[147] = 8'd241; M[148] = 8'd16; M[149] = 8'd232; M[150] = 8'd194; M[151] = 8'd201; 
M[208] = 8'd191; M[209] = 8'd186; M[210] = 8'd199; M[211] = 8'd250; M[212] = 8'd26; M[213] = 8'd234; M[214] = 8'd198; M[215] = 8'd197; 
M[272] = 8'd195; M[273] = 8'd189; M[274] = 8'd196; M[275] = 8'd232; M[276] = 8'd254; M[277] = 8'd216; M[278] = 8'd196; M[279] = 8'd198; 
M[336] = 8'd207; M[337] = 8'd193; M[338] = 8'd188; M[339] = 8'd198; M[340] = 8'd205; M[341] = 8'd196; M[342] = 8'd186; M[343] = 8'd203; 
M[400] = 8'd213; M[401] = 8'd199; M[402] = 8'd192; M[403] = 8'd187; M[404] = 8'd183; M[405] = 8'd189; M[406] = 8'd193; M[407] = 8'd211; 
M[464] = 8'd215; M[465] = 8'd207; M[466] = 8'd197; M[467] = 8'd196; M[468] = 8'd193; M[469] = 8'd204; M[470] = 8'd206; M[471] = 8'd222; 

M[24] = 8'd180; M[25] = 8'd183; M[26] = 8'd189; M[27] = 8'd194; M[28] = 8'd198; M[29] = 8'd189; M[30] = 8'd192; M[31] = 8'd201; 
M[88] = 8'd191; M[89] = 8'd187; M[90] = 8'd183; M[91] = 8'd218; M[92] = 8'd237; M[93] = 8'd213; M[94] = 8'd197; M[95] = 8'd200; 
M[152] = 8'd190; M[153] = 8'd187; M[154] = 8'd196; M[155] = 8'd241; M[156] = 8'd16; M[157] = 8'd232; M[158] = 8'd194; M[159] = 8'd201; 
M[216] = 8'd191; M[217] = 8'd186; M[218] = 8'd199; M[219] = 8'd250; M[220] = 8'd26; M[221] = 8'd234; M[222] = 8'd198; M[223] = 8'd197; 
M[280] = 8'd195; M[281] = 8'd189; M[282] = 8'd196; M[283] = 8'd232; M[284] = 8'd254; M[285] = 8'd216; M[286] = 8'd196; M[287] = 8'd198; 
M[344] = 8'd207; M[345] = 8'd193; M[346] = 8'd188; M[347] = 8'd198; M[348] = 8'd205; M[349] = 8'd196; M[350] = 8'd186; M[351] = 8'd203; 
M[408] = 8'd213; M[409] = 8'd199; M[410] = 8'd192; M[411] = 8'd187; M[412] = 8'd183; M[413] = 8'd189; M[414] = 8'd193; M[415] = 8'd211; 
M[472] = 8'd215; M[473] = 8'd207; M[474] = 8'd197; M[475] = 8'd196; M[476] = 8'd193; M[477] = 8'd204; M[478] = 8'd206; M[479] = 8'd222; 

M[32] = 8'd180; M[33] = 8'd183; M[34] = 8'd189; M[35] = 8'd194; M[36] = 8'd198; M[37] = 8'd189; M[38] = 8'd192; M[39] = 8'd201; 
M[96] = 8'd191; M[97] = 8'd187; M[98] = 8'd183; M[99] = 8'd218; M[100] = 8'd237; M[101] = 8'd213; M[102] = 8'd197; M[103] = 8'd200; 
M[160] = 8'd190; M[161] = 8'd187; M[162] = 8'd196; M[163] = 8'd241; M[164] = 8'd16; M[165] = 8'd232; M[166] = 8'd194; M[167] = 8'd201; 
M[224] = 8'd191; M[225] = 8'd186; M[226] = 8'd199; M[227] = 8'd250; M[228] = 8'd26; M[229] = 8'd234; M[230] = 8'd198; M[231] = 8'd197; 
M[288] = 8'd195; M[289] = 8'd189; M[290] = 8'd196; M[291] = 8'd232; M[292] = 8'd254; M[293] = 8'd216; M[294] = 8'd196; M[295] = 8'd198; 
M[352] = 8'd207; M[353] = 8'd193; M[354] = 8'd188; M[355] = 8'd198; M[356] = 8'd205; M[357] = 8'd196; M[358] = 8'd186; M[359] = 8'd203; 
M[416] = 8'd213; M[417] = 8'd199; M[418] = 8'd192; M[419] = 8'd187; M[420] = 8'd183; M[421] = 8'd189; M[422] = 8'd193; M[423] = 8'd211; 
M[480] = 8'd215; M[481] = 8'd207; M[482] = 8'd197; M[483] = 8'd196; M[484] = 8'd193; M[485] = 8'd204; M[486] = 8'd206; M[487] = 8'd222; 

M[40] = 8'd180; M[41] = 8'd183; M[42] = 8'd189; M[43] = 8'd194; M[44] = 8'd198; M[45] = 8'd189; M[46] = 8'd192; M[47] = 8'd201; 
M[104] = 8'd191; M[105] = 8'd187; M[106] = 8'd183; M[107] = 8'd218; M[108] = 8'd237; M[109] = 8'd213; M[110] = 8'd197; M[111] = 8'd200; 
M[168] = 8'd190; M[169] = 8'd187; M[170] = 8'd196; M[171] = 8'd241; M[172] = 8'd16; M[173] = 8'd232; M[174] = 8'd194; M[175] = 8'd201; 
M[232] = 8'd191; M[233] = 8'd186; M[234] = 8'd199; M[235] = 8'd250; M[236] = 8'd26; M[237] = 8'd234; M[238] = 8'd198; M[239] = 8'd197; 
M[296] = 8'd195; M[297] = 8'd189; M[298] = 8'd196; M[299] = 8'd232; M[300] = 8'd254; M[301] = 8'd216; M[302] = 8'd196; M[303] = 8'd198; 
M[360] = 8'd207; M[361] = 8'd193; M[362] = 8'd188; M[363] = 8'd198; M[364] = 8'd205; M[365] = 8'd196; M[366] = 8'd186; M[367] = 8'd203; 
M[424] = 8'd213; M[425] = 8'd199; M[426] = 8'd192; M[427] = 8'd187; M[428] = 8'd183; M[429] = 8'd189; M[430] = 8'd193; M[431] = 8'd211; 
M[488] = 8'd215; M[489] = 8'd207; M[490] = 8'd197; M[491] = 8'd196; M[492] = 8'd193; M[493] = 8'd204; M[494] = 8'd206; M[495] = 8'd222; 

M[48] = 8'd180; M[49] = 8'd183; M[50] = 8'd189; M[51] = 8'd194; M[52] = 8'd198; M[53] = 8'd189; M[54] = 8'd192; M[55] = 8'd201; 
M[112] = 8'd191; M[113] = 8'd187; M[114] = 8'd183; M[115] = 8'd218; M[116] = 8'd237; M[117] = 8'd213; M[118] = 8'd197; M[119] = 8'd200; 
M[176] = 8'd190; M[177] = 8'd187; M[178] = 8'd196; M[179] = 8'd241; M[180] = 8'd16; M[181] = 8'd232; M[182] = 8'd194; M[183] = 8'd201; 
M[240] = 8'd191; M[241] = 8'd186; M[242] = 8'd199; M[243] = 8'd250; M[244] = 8'd26; M[245] = 8'd234; M[246] = 8'd198; M[247] = 8'd197; 
M[304] = 8'd195; M[305] = 8'd189; M[306] = 8'd196; M[307] = 8'd232; M[308] = 8'd254; M[309] = 8'd216; M[310] = 8'd196; M[311] = 8'd198; 
M[368] = 8'd207; M[369] = 8'd193; M[370] = 8'd188; M[371] = 8'd198; M[372] = 8'd205; M[373] = 8'd196; M[374] = 8'd186; M[375] = 8'd203; 
M[432] = 8'd213; M[433] = 8'd199; M[434] = 8'd192; M[435] = 8'd187; M[436] = 8'd183; M[437] = 8'd189; M[438] = 8'd193; M[439] = 8'd211; 
M[496] = 8'd215; M[497] = 8'd207; M[498] = 8'd197; M[499] = 8'd196; M[500] = 8'd193; M[501] = 8'd204; M[502] = 8'd206; M[503] = 8'd222; 

M[56] = 8'd180; M[57] = 8'd183; M[58] = 8'd189; M[59] = 8'd194; M[60] = 8'd198; M[61] = 8'd189; M[62] = 8'd192; M[63] = 8'd201; 
M[120] = 8'd191; M[121] = 8'd187; M[122] = 8'd183; M[123] = 8'd218; M[124] = 8'd237; M[125] = 8'd213; M[126] = 8'd197; M[127] = 8'd200; 
M[184] = 8'd190; M[185] = 8'd187; M[186] = 8'd196; M[187] = 8'd241; M[188] = 8'd16; M[189] = 8'd232; M[190] = 8'd194; M[191] = 8'd201; 
M[248] = 8'd191; M[249] = 8'd186; M[250] = 8'd199; M[251] = 8'd250; M[252] = 8'd26; M[253] = 8'd234; M[254] = 8'd198; M[255] = 8'd197; 
M[312] = 8'd195; M[313] = 8'd189; M[314] = 8'd196; M[315] = 8'd232; M[316] = 8'd254; M[317] = 8'd216; M[318] = 8'd196; M[319] = 8'd198; 
M[376] = 8'd207; M[377] = 8'd193; M[378] = 8'd188; M[379] = 8'd198; M[380] = 8'd205; M[381] = 8'd196; M[382] = 8'd186; M[383] = 8'd203; 
M[440] = 8'd213; M[441] = 8'd199; M[442] = 8'd192; M[443] = 8'd187; M[444] = 8'd183; M[445] = 8'd189; M[446] = 8'd193; M[447] = 8'd211; 
M[504] = 8'd215; M[505] = 8'd207; M[506] = 8'd197; M[507] = 8'd196; M[508] = 8'd193; M[509] = 8'd204; M[510] = 8'd206; M[511] = 8'd222;
//I[1] = M[0];
rst[1:Total_MCUs] = {Total_MCUs{1'b1}};
//rst[2] = 1'b1;
//rst[3] = 1'b1;
//O=2432'd0;
en[1:Total_MCUs] = {1'b1,{Total_MCUs-1{1'b0}}};
//en[2] = 1'b0;
//en[3] = 1'b0;
dc_in[1] = 14'd0;
MCU_ctr = 11'd0;
first_MCU = 1'b1;
change = 1'b1;
start = 1'b0;
st = 1'b0;
start_MCU[1:Total_MCUs] = {Total_MCUs{1'b0}};
//start_MCU[2] = 1'b0;
//start_MCU[3] = 1'b0;
end

always begin
#1 clk=~clk;
//always@(negedge clk)
//rst=0;
//I = M[0];
end

always@(posedge clk) begin
// defaults
//    I1 <= I1;
//    I2 <= I2;
    
//    en1 <= 1'b0;
//    en2 <= 1'b0;
    if(start == 1'b0) begin
        start <= 1'b1;
        present_MCU <= 10'd1;
        en[1] <= 1'b1;
        I[1] <= M[0];           //Input is supplied as soon as enable is 1
//        overall_ctr <= 20'd1;
        rst[1:Total_MCUs] <= {Total_MCUs{1'b0}};
//        rst[2] <= 1'b0;
//        rst[3] <= 1'b0;
        start_MCU[1] <= 1'b1;
    end

    if(start == 1'b1) begin
        overall_ctr = overall_ctr + 1'b1; 
    end

    st <= start;    // Helpful to decide transition
    
    if(overall_ctr[2:0] == 3'b000 && st == 1) begin
        if(present_MCU == Total_MCUs) begin  // last MCU
            present_MCU = 10'd1;    //<
            I[1] = M[overall_ctr];
            en[Total_MCUs] = 1'b0;  // enables
            en[1] = 1'b1;
            first_MCU = 1'b1;
        end
        else begin                      // MCU 1-> MCU 2, 2->3
            present_MCU = present_MCU + 1'b1;//<
            I[present_MCU] = M[overall_ctr];
            en[present_MCU] = 1'b1;
            en[present_MCU - 1] = 1'b0;
            first_MCU = 1'b0;//<
            start_MCU[present_MCU] <= 1'b1;// + 1
        end
    end
    else begin
            I[present_MCU] = M[overall_ctr];
            en[present_MCU] = 1'b1;
    end
end



always@(posedge(Valid_output[1])) begin
    dc_in[2] <= dc_out[1];
end

always@(posedge(Valid_output[2])) begin
    dc_in[3] <= dc_out[2];
end


DCT_2D MCU_1(I[1], rst[1], clk, en[1], dc_in[1], start_MCU[1], ready[1], O[1], done[1], dc_out[1], first_MCU, Valid_output[1]);
DCT_2D MCU_2(I[2], rst[2], clk, en[2], dc_in[2], start_MCU[2], ready[2], O[2], done[2], dc_out[2], first_MCU, Valid_output[2]);
DCT_2D MCU_3(I[3], rst[3], clk, en[3], dc_in[3], start_MCU[3], ready[3], O[3], done[3], dc_out[3], first_MCU, Valid_output[3]);
DCT_2D MCU_4(I[4], rst[4], clk, en[4], dc_in[4], start_MCU[4], ready[4], O[4], done[4], dc_out[4], first_MCU, Valid_output[4]);
DCT_2D MCU_5(I[5], rst[5], clk, en[5], dc_in[5], start_MCU[5], ready[5], O[5], done[5], dc_out[5], first_MCU, Valid_output[5]);
DCT_2D MCU_6(I[6], rst[6], clk, en[6], dc_in[6], start_MCU[6], ready[6], O[6], done[6], dc_out[6], first_MCU, Valid_output[6]);
DCT_2D MCU_7(I[7], rst[7], clk, en[7], dc_in[7], start_MCU[7], ready[7], O[7], done[7], dc_out[7], first_MCU, Valid_output[7]);
DCT_2D MCU_8(I[8], rst[8], clk, en[8], dc_in[8], start_MCU[8], ready[8], O[8], done[8], dc_out[8], first_MCU, Valid_output[8]);
endmodule
