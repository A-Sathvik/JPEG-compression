`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.04.2021 14:07:32
// Design Name: 
// Module Name: Huffman_encoding
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// OM
//////////////////////////////////////////////////////////////////////////////////


module Huffman_encoding(clk,dc,dc_value,run,Size,Suffix_code,final_term,After_H);
input clk,dc;   // Signal dc conveys whether the Coefficient is dc or not(i.e, ac)
input [7:0] dc_value;
input [3:0] run;      // for example 0 in (0,15)
input [2:0] Size;     // size of suffix code of 15
input [6:0] Suffix_code;    // Code for 15
input final_term;
output reg [0:22] After_H;    // huffman encoded bit string
always@(posedge clk) begin
if(final_term == 1'b1) begin
    After_H <= {4'b1010,19'd0};
end
else begin
    if(dc == 1'b1) begin
        case(dc_value)
            8'd192: After_H <= {12'b111100111111, 11'd0}; // -64
            8'd193: After_H <= {10'b1110000000, 13'd0}; // -63
            8'd194: After_H <= {10'b1110000001, 13'd0}; // -62
            8'd195: After_H <= {10'b1110000010, 13'd0}; // -61
            8'd196: After_H <= {10'b1110000011, 13'd0}; // -60
            8'd197: After_H <= {10'b1110000100, 13'd0}; // -59
            8'd198: After_H <= {10'b1110000101, 13'd0}; // -58
            8'd199: After_H <= {10'b1110000110, 13'd0}; // -57
            8'd200: After_H <= {10'b1110000111, 13'd0}; // -56
            8'd201: After_H <= {10'b1110001000, 13'd0}; // -55
            8'd202: After_H <= {10'b1110001001, 13'd0}; // -54
            8'd203: After_H <= {10'b1110001010, 13'd0}; // -53
            8'd204: After_H <= {10'b1110001011, 13'd0}; // -52
            8'd205: After_H <= {10'b1110001100, 13'd0}; // -51
            8'd206: After_H <= {10'b1110001101, 13'd0}; // -50
            8'd207: After_H <= {10'b1110001110, 13'd0}; // -49
            8'd208: After_H <= {10'b1110001111, 13'd0}; // -48
            8'd209: After_H <= {10'b1110010000, 13'd0}; // -47
            8'd210: After_H <= {10'b1110010001, 13'd0}; // -46
            8'd211: After_H <= {10'b1110010010, 13'd0}; // -45
            8'd212: After_H <= {10'b1110010011, 13'd0}; // -44
            8'd213: After_H <= {10'b1110010100, 13'd0}; // -43
            8'd214: After_H <= {10'b1110010101, 13'd0}; // -42
            8'd215: After_H <= {10'b1110010110, 13'd0}; // -41
            8'd216: After_H <= {10'b1110010111, 13'd0}; // -40
            8'd217: After_H <= {10'b1110011000, 13'd0}; // -39
            8'd218: After_H <= {10'b1110011001, 13'd0}; // -38
            8'd219: After_H <= {10'b1110011010, 13'd0}; // -37
            8'd220: After_H <= {10'b1110011011, 13'd0}; // -36
            8'd221: After_H <= {10'b1110011100, 13'd0}; // -35
            8'd222: After_H <= {10'b1110011101, 13'd0}; // -34
            8'd223: After_H <= {10'b1110011110, 13'd0}; // -33
            8'd224: After_H <= {10'b1110011111, 13'd0}; // -32
            8'd225: After_H <= {8'b11000000, 15'd0}; // -31
            8'd226: After_H <= {8'b11000001, 15'd0}; // -30
            8'd227: After_H <= {8'b11000010, 15'd0}; // -29
            8'd228: After_H <= {8'b11000011, 15'd0}; // -28
            8'd229: After_H <= {8'b11000100, 15'd0}; // -27
            8'd230: After_H <= {8'b11000101, 15'd0}; // -26
            8'd231: After_H <= {8'b11000110, 15'd0}; // -25
            8'd232: After_H <= {8'b11000111, 15'd0}; // -24
            8'd233: After_H <= {8'b11001000, 15'd0}; // -23
            8'd234: After_H <= {8'b11001001, 15'd0}; // -22
            8'd235: After_H <= {8'b11001010, 15'd0}; // -21
            8'd236: After_H <= {8'b11001011, 15'd0}; // -20
            8'd237: After_H <= {8'b11001100, 15'd0}; // -19
            8'd238: After_H <= {8'b11001101, 15'd0}; // -18
            8'd239: After_H <= {8'b11001110, 15'd0}; // -17
            8'd240: After_H <= {8'b11001111, 15'd0}; // -16
            8'd241: After_H <= {7'b1010000, 16'd0}; // -15
            8'd242: After_H <= {7'b1010001, 16'd0}; // -14
            8'd243: After_H <= {7'b1010010, 16'd0}; // -13
            8'd244: After_H <= {7'b1010011, 16'd0}; // -12
            8'd245: After_H <= {7'b1010100, 16'd0}; // -11
            8'd246: After_H <= {7'b1010101, 16'd0}; // -10
            8'd247: After_H <= {7'b1010110, 16'd0}; // -9
            8'd248: After_H <= {7'b1010111, 16'd0}; // -8
            8'd249: After_H <= {6'b100000, 17'd0}; // -7
            8'd250: After_H <= {6'b100001, 17'd0}; // -6
            8'd251: After_H <= {6'b100010, 17'd0}; // -5
            8'd252: After_H <= {6'b100011, 17'd0}; // -4
            8'd253: After_H <= {5'b01100, 18'd0}; // -3
            8'd254: After_H <= {5'b01101, 18'd0}; // -2
            8'd255: After_H <= {4'b0100, 19'd0}; // -1
            8'd0: After_H <= {2'b00, 21'd0}; // 0
            8'd1: After_H <= {4'b0101, 19'd0}; // 1
            8'd2: After_H <= {5'b01110, 18'd0}; // 2
            8'd3: After_H <= {5'b01111, 18'd0}; // 3
            8'd4: After_H <= {6'b100100, 17'd0}; // 4
            8'd5: After_H <= {6'b100101, 17'd0}; // 5
            8'd6: After_H <= {6'b100110, 17'd0}; // 6
            8'd7: After_H <= {6'b100111, 17'd0}; // 7
            8'd8: After_H <= {7'b1011000, 16'd0}; // 8
            8'd9: After_H <= {7'b1011001, 16'd0}; // 9
            8'd10: After_H <= {7'b1011010, 16'd0}; // 10
            8'd11: After_H <= {7'b1011011, 16'd0}; // 11
            8'd12: After_H <= {7'b1011100, 16'd0}; // 12
            8'd13: After_H <= {7'b1011101, 16'd0}; // 13
            8'd14: After_H <= {7'b1011110, 16'd0}; // 14
            8'd15: After_H <= {7'b1011111, 16'd0}; // 15
            8'd16: After_H <= {8'b11010000, 15'd0}; // 16
            8'd17: After_H <= {8'b11010001, 15'd0}; // 17
            8'd18: After_H <= {8'b11010010, 15'd0}; // 18
            8'd19: After_H <= {8'b11010011, 15'd0}; // 19
            8'd20: After_H <= {8'b11010100, 15'd0}; // 20
            8'd21: After_H <= {8'b11010101, 15'd0}; // 21
            8'd22: After_H <= {8'b11010110, 15'd0}; // 22
            8'd23: After_H <= {8'b11010111, 15'd0}; // 23
            8'd24: After_H <= {8'b11011000, 15'd0}; // 24
            8'd25: After_H <= {8'b11011001, 15'd0}; // 25
            8'd26: After_H <= {8'b11011010, 15'd0}; // 26
            8'd27: After_H <= {8'b11011011, 15'd0}; // 27
            8'd28: After_H <= {8'b11011100, 15'd0}; // 28
            8'd29: After_H <= {8'b11011101, 15'd0}; // 29
            8'd30: After_H <= {8'b11011110, 15'd0}; // 30
            8'd31: After_H <= {8'b11011111, 15'd0}; // 31
            8'd32: After_H <= {10'b1110100000, 13'd0}; // 32
            8'd33: After_H <= {10'b1110100001, 13'd0}; // 33
            8'd34: After_H <= {10'b1110100010, 13'd0}; // 34
            8'd35: After_H <= {10'b1110100011, 13'd0}; // 35
            8'd36: After_H <= {10'b1110100100, 13'd0}; // 36
            8'd37: After_H <= {10'b1110100101, 13'd0}; // 37
            8'd38: After_H <= {10'b1110100110, 13'd0}; // 38
            8'd39: After_H <= {10'b1110100111, 13'd0}; // 39
            8'd40: After_H <= {10'b1110101000, 13'd0}; // 40
            8'd41: After_H <= {10'b1110101001, 13'd0}; // 41
            8'd42: After_H <= {10'b1110101010, 13'd0}; // 42
            8'd43: After_H <= {10'b1110101011, 13'd0}; // 43
            8'd44: After_H <= {10'b1110101100, 13'd0}; // 44
            8'd45: After_H <= {10'b1110101101, 13'd0}; // 45
            8'd46: After_H <= {10'b1110101110, 13'd0}; // 46
            8'd47: After_H <= {10'b1110101111, 13'd0}; // 47
            8'd48: After_H <= {10'b1110110000, 13'd0}; // 48
            8'd49: After_H <= {10'b1110110001, 13'd0}; // 49
            8'd50: After_H <= {10'b1110110010, 13'd0}; // 50
            8'd51: After_H <= {10'b1110110011, 13'd0}; // 51
            8'd52: After_H <= {10'b1110110100, 13'd0}; // 52
            8'd53: After_H <= {10'b1110110101, 13'd0}; // 53
            8'd54: After_H <= {10'b1110110110, 13'd0}; // 54
            8'd55: After_H <= {10'b1110110111, 13'd0}; // 55
            8'd56: After_H <= {10'b1110111000, 13'd0}; // 56
            8'd57: After_H <= {10'b1110111001, 13'd0}; // 57
            8'd58: After_H <= {10'b1110111010, 13'd0}; // 58
            8'd59: After_H <= {10'b1110111011, 13'd0}; // 59
            8'd60: After_H <= {10'b1110111100, 13'd0}; // 60
            8'd61: After_H <= {10'b1110111101, 13'd0}; // 61
            8'd62: After_H <= {10'b1110111110, 13'd0}; // 62
            8'd63: After_H <= {10'b1110111111, 13'd0}; // 63
            default : After_H <= {23{1'b0}};
        endcase
    end
    else begin  // For ac values
        case ({run,Size})
        {4'b0000,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 0/0
        {4'b0000,3'b001}: After_H <= {2'b00, Suffix_code[0], 20'd0}; // 0/1
        {4'b0000,3'b010}: After_H <= {2'b01, Suffix_code[1:0], 19'd0}; // 0/2
        {4'b0000,3'b011}: After_H <= {3'b100, Suffix_code[2:0], 17'd0}; // 0/3
        {4'b0000,3'b100}: After_H <= {4'b1011, Suffix_code[3:0], 15'd0}; // 0/4
        {4'b0000,3'b101}: After_H <= {5'b11010, Suffix_code[4:0], 13'd0}; // 0/5
        {4'b0000,3'b110}: After_H <= {7'b1111000, Suffix_code[5:0], 10'd0}; // 0/6
        {4'b0000,3'b111}: After_H <= {8'b11111000, Suffix_code[6:0], 8'd0}; // 0/7
        {4'b0001,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 1/0
        {4'b0001,3'b001}: After_H <= {4'b1100, Suffix_code[0], 18'd0}; // 1/1
        {4'b0001,3'b010}: After_H <= {5'b11011, Suffix_code[1:0], 16'd0}; // 1/2
        {4'b0001,3'b011}: After_H <= {7'b1111001, Suffix_code[2:0], 13'd0}; // 1/3
        {4'b0001,3'b100}: After_H <= {9'b111110110, Suffix_code[3:0], 10'd0}; // 1/4
        {4'b0001,3'b101}: After_H <= {11'b11111110110, Suffix_code[4:0], 7'd0}; // 1/5
        {4'b0001,3'b110}: After_H <= {16'b1111111110000100, Suffix_code[5:0], 1'd0}; // 1/6
        {4'b0001,3'b111}: After_H <= {16'b1111111110000101, Suffix_code[6:0]}; // 1/7
        {4'b0010,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 2/0
        {4'b0010,3'b001}: After_H <= {5'b11100, Suffix_code[0], 17'd0}; // 2/1
        {4'b0010,3'b010}: After_H <= {8'b11111001, Suffix_code[1:0], 13'd0}; // 2/2
        {4'b0010,3'b011}: After_H <= {10'b1111110111, Suffix_code[2:0], 10'd0}; // 2/3
        {4'b0010,3'b100}: After_H <= {12'b111111110100, Suffix_code[3:0], 7'd0}; // 2/4
        {4'b0010,3'b101}: After_H <= {16'b1111111110001001, Suffix_code[4:0], 2'd0}; // 2/5
        {4'b0010,3'b110}: After_H <= {16'b1111111110001010, Suffix_code[5:0], 1'd0}; // 2/6
        {4'b0010,3'b111}: After_H <= {16'b1111111110001011, Suffix_code[6:0]}; // 2/7
        {4'b0011,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 3/0
        {4'b0011,3'b001}: After_H <= {6'b111010, Suffix_code[0], 16'd0}; // 3/1
        {4'b0011,3'b010}: After_H <= {9'b111110111, Suffix_code[1:0], 12'd0}; // 3/2
        {4'b0011,3'b011}: After_H <= {12'b111111110101, Suffix_code[2:0], 8'd0}; // 3/3
        {4'b0011,3'b100}: After_H <= {16'b1111111110001111, Suffix_code[3:0], 3'd0}; // 3/4
        {4'b0011,3'b101}: After_H <= {16'b1111111110010000, Suffix_code[4:0], 2'd0}; // 3/5
        {4'b0011,3'b110}: After_H <= {16'b1111111110010001, Suffix_code[5:0], 1'd0}; // 3/6
        {4'b0011,3'b111}: After_H <= {16'b1111111110010010, Suffix_code[6:0]}; // 3/7
        {4'b0100,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 4/0
        {4'b0100,3'b001}: After_H <= {6'b111011, Suffix_code[0], 16'd0}; // 4/1
        {4'b0100,3'b010}: After_H <= {10'b1111111000, Suffix_code[1:0], 11'd0}; // 4/2
        {4'b0100,3'b011}: After_H <= {16'b1111111110010110, Suffix_code[2:0], 4'd0}; // 4/3
        {4'b0100,3'b100}: After_H <= {16'b1111111110010111, Suffix_code[3:0], 3'd0}; // 4/4
        {4'b0100,3'b101}: After_H <= {16'b1111111110011000, Suffix_code[4:0], 2'd0}; // 4/5
        {4'b0100,3'b110}: After_H <= {16'b1111111110011001, Suffix_code[5:0], 1'd0}; // 4/6
        {4'b0100,3'b111}: After_H <= {16'b1111111110011010, Suffix_code[6:0]}; // 4/7
        {4'b0101,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 5/0
        {4'b0101,3'b001}: After_H <= {7'b1111010, Suffix_code[0], 15'd0}; // 5/1
        {4'b0101,3'b010}: After_H <= {11'b11111110111, Suffix_code[1:0], 10'd0}; // 5/2
        {4'b0101,3'b011}: After_H <= {16'b1111111110011110, Suffix_code[2:0], 4'd0}; // 5/3
        {4'b0101,3'b100}: After_H <= {16'b1111111110011111, Suffix_code[3:0], 3'd0}; // 5/4
        {4'b0101,3'b101}: After_H <= {16'b1111111110100000, Suffix_code[4:0], 2'd0}; // 5/5
        {4'b0101,3'b110}: After_H <= {16'b1111111110100001, Suffix_code[5:0], 1'd0}; // 5/6
        {4'b0101,3'b111}: After_H <= {16'b1111111110100010, Suffix_code[6:0]}; // 5/7
        {4'b0110,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 6/0
        {4'b0110,3'b001}: After_H <= {7'b1111011, Suffix_code[0], 15'd0}; // 6/1
        {4'b0110,3'b010}: After_H <= {12'b111111110110, Suffix_code[1:0], 9'd0}; // 6/2
        {4'b0110,3'b011}: After_H <= {16'b1111111110100110, Suffix_code[2:0], 4'd0}; // 6/3
        {4'b0110,3'b100}: After_H <= {16'b1111111110100111, Suffix_code[3:0], 3'd0}; // 6/4
        {4'b0110,3'b101}: After_H <= {16'b1111111110101000, Suffix_code[4:0], 2'd0}; // 6/5
        {4'b0110,3'b110}: After_H <= {16'b1111111110101001, Suffix_code[5:0], 1'd0}; // 6/6
        {4'b0110,3'b111}: After_H <= {16'b1111111110101010, Suffix_code[6:0]}; // 6/7
        {4'b0111,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 7/0
        {4'b0111,3'b001}: After_H <= {8'b11111010, Suffix_code[0], 14'd0}; // 7/1
        {4'b0111,3'b010}: After_H <= {12'b111111110111, Suffix_code[1:0], 9'd0}; // 7/2
        {4'b0111,3'b011}: After_H <= {16'b1111111110101110, Suffix_code[2:0], 4'd0}; // 7/3
        {4'b0111,3'b100}: After_H <= {16'b1111111110101111, Suffix_code[3:0], 3'd0}; // 7/4
        {4'b0111,3'b101}: After_H <= {16'b1111111110110000, Suffix_code[4:0], 2'd0}; // 7/5
        {4'b0111,3'b110}: After_H <= {16'b1111111110110001, Suffix_code[5:0], 1'd0}; // 7/6
        {4'b0111,3'b111}: After_H <= {16'b1111111110110010, Suffix_code[6:0]}; // 7/7
        {4'b1000,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 8/0
        {4'b1000,3'b001}: After_H <= {9'b111111000, Suffix_code[0], 13'd0}; // 8/1
        {4'b1000,3'b010}: After_H <= {15'b111111111000000, Suffix_code[1:0], 6'd0}; // 8/2
        {4'b1000,3'b011}: After_H <= {16'b1111111110110110, Suffix_code[2:0], 4'd0}; // 8/3
        {4'b1000,3'b100}: After_H <= {16'b1111111110110111, Suffix_code[3:0], 3'd0}; // 8/4
        {4'b1000,3'b101}: After_H <= {16'b1111111110111000, Suffix_code[4:0], 2'd0}; // 8/5
        {4'b1000,3'b110}: After_H <= {16'b1111111110111001, Suffix_code[5:0], 1'd0}; // 8/6
        {4'b1000,3'b111}: After_H <= {16'b1111111110111010, Suffix_code[6:0]}; // 8/7
        {4'b1001,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 9/0
        {4'b1001,3'b001}: After_H <= {9'b111111001, Suffix_code[0], 13'd0}; // 9/1
        {4'b1001,3'b010}: After_H <= {16'b1111111110111110, Suffix_code[1:0], 5'd0}; // 9/2
        {4'b1001,3'b011}: After_H <= {16'b1111111110111111, Suffix_code[2:0], 4'd0}; // 9/3
        {4'b1001,3'b100}: After_H <= {16'b1111111111000000, Suffix_code[3:0], 3'd0}; // 9/4
        {4'b1001,3'b101}: After_H <= {16'b1111111111000001, Suffix_code[4:0], 2'd0}; // 9/5
        {4'b1001,3'b110}: After_H <= {16'b1111111111000010, Suffix_code[5:0], 1'd0}; // 9/6
        {4'b1001,3'b111}: After_H <= {16'b1111111111000011, Suffix_code[6:0]}; // 9/7
        {4'b1010,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 10/0
        {4'b1010,3'b001}: After_H <= {9'b111111010, Suffix_code[0], 13'd0}; // 10/1
        {4'b1010,3'b010}: After_H <= {16'b1111111111000111, Suffix_code[1:0], 5'd0}; // 10/2
        {4'b1010,3'b011}: After_H <= {16'b1111111111001000, Suffix_code[2:0], 4'd0}; // 10/3
        {4'b1010,3'b100}: After_H <= {16'b1111111111001001, Suffix_code[3:0], 3'd0}; // 10/4
        {4'b1010,3'b101}: After_H <= {16'b1111111111001010, Suffix_code[4:0], 2'd0}; // 10/5
        {4'b1010,3'b110}: After_H <= {16'b1111111111001011, Suffix_code[5:0], 1'd0}; // 10/6
        {4'b1010,3'b111}: After_H <= {16'b1111111111001100, Suffix_code[6:0]}; // 10/7
        {4'b1011,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 11/0
        {4'b1011,3'b001}: After_H <= {10'b1111111001, Suffix_code[0], 12'd0}; // 11/1
        {4'b1011,3'b010}: After_H <= {16'b1111111111010000, Suffix_code[1:0], 5'd0}; // 11/2
        {4'b1011,3'b011}: After_H <= {16'b1111111111010001, Suffix_code[2:0], 4'd0}; // 11/3
        {4'b1011,3'b100}: After_H <= {16'b1111111111010010, Suffix_code[3:0], 3'd0}; // 11/4
        {4'b1011,3'b101}: After_H <= {16'b1111111111010011, Suffix_code[4:0], 2'd0}; // 11/5
        {4'b1011,3'b110}: After_H <= {16'b1111111111010100, Suffix_code[5:0], 1'd0}; // 11/6
        {4'b1011,3'b111}: After_H <= {16'b1111111111010101, Suffix_code[6:0]}; // 11/7
        {4'b1100,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 12/0
        {4'b1100,3'b001}: After_H <= {10'b1111111010, Suffix_code[0], 12'd0}; // 12/1
        {4'b1100,3'b010}: After_H <= {16'b1111111111011001, Suffix_code[1:0], 5'd0}; // 12/2
        {4'b1100,3'b011}: After_H <= {16'b1111111111011010, Suffix_code[2:0], 4'd0}; // 12/3
        {4'b1100,3'b100}: After_H <= {16'b1111111111011011, Suffix_code[3:0], 3'd0}; // 12/4
        {4'b1100,3'b101}: After_H <= {16'b1111111111011100, Suffix_code[4:0], 2'd0}; // 12/5
        {4'b1100,3'b110}: After_H <= {16'b1111111111011101, Suffix_code[5:0], 1'd0}; // 12/6
        {4'b1100,3'b111}: After_H <= {16'b1111111111011110, Suffix_code[6:0]}; // 12/7
        {4'b1101,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 13/0
        {4'b1101,3'b001}: After_H <= {11'b11111111000, Suffix_code[0], 11'd0}; // 13/1
        {4'b1101,3'b010}: After_H <= {16'b1111111111100010, Suffix_code[1:0], 5'd0}; // 13/2
        {4'b1101,3'b011}: After_H <= {16'b1111111111100011, Suffix_code[2:0], 4'd0}; // 13/3
        {4'b1101,3'b100}: After_H <= {16'b1111111111100100, Suffix_code[3:0], 3'd0}; // 13/4
        {4'b1101,3'b101}: After_H <= {16'b1111111111100101, Suffix_code[4:0], 2'd0}; // 13/5
        {4'b1101,3'b110}: After_H <= {16'b1111111111100110, Suffix_code[5:0], 1'd0}; // 13/6
        {4'b1101,3'b111}: After_H <= {16'b1111111111100111, Suffix_code[6:0]}; // 13/7
        {4'b1110,3'b000}: After_H <= {4'b1010, 19'd0};  // End of input 14/0
        {4'b1110,3'b001}: After_H <= {16'b1111111111101011, Suffix_code[0], 6'd0}; // 14/1
        {4'b1110,3'b010}: After_H <= {16'b1111111111101100, Suffix_code[1:0], 5'd0}; // 14/2
        {4'b1110,3'b011}: After_H <= {16'b1111111111101101, Suffix_code[2:0], 4'd0}; // 14/3
        {4'b1110,3'b100}: After_H <= {16'b1111111111101110, Suffix_code[3:0], 3'd0}; // 14/4
        {4'b1110,3'b101}: After_H <= {16'b1111111111101111, Suffix_code[4:0], 2'd0}; // 14/5
        {4'b1110,3'b110}: After_H <= {16'b1111111111110000, Suffix_code[5:0], 1'd0}; // 14/6
        {4'b1110,3'b111}: After_H <= {16'b1111111111110001, Suffix_code[6:0]}; // 14/7
        {4'b1111,3'b000}: After_H <= {11'b11111111001,12'd0}; // 15/0
        {4'b1111,3'b001}: After_H <= {16'b1111111111110101, Suffix_code[0], 6'd0}; // 15/1
        {4'b1111,3'b010}: After_H <= {16'b1111111111110110, Suffix_code[1:0], 5'd0}; // 15/2
        {4'b1111,3'b011}: After_H <= {16'b1111111111110111, Suffix_code[2:0], 4'd0}; // 15/3
        {4'b1111,3'b100}: After_H <= {16'b1111111111111000, Suffix_code[3:0], 3'd0}; // 15/4
        {4'b1111,3'b101}: After_H <= {16'b1111111111111001, Suffix_code[4:0], 2'd0}; // 15/5
        {4'b1111,3'b110}: After_H <= {16'b1111111111111010, Suffix_code[5:0], 1'd0}; // 15/6
        {4'b1111,3'b111}: After_H <= {16'b111111111111101, Suffix_code[6:0]}; // 15/7
        endcase
    end // A.C terms loop
end // final_term, else loop
end
endmodule
